-- #################################################################################################
-- # << NEORV32 for the iCEBreaker FPGA Board >>                                                   #
-- # ********************************************************************************************* #
-- # FPGA:  Lattice iCE40UP5k                                                                      #
-- # Board: https://github.com/icebreaker-fpga/icebreaker                                          #
-- # ********************************************************************************************* #
-- # BSD 3-Clause License                                                                          #
-- #                                                                                               #
-- # The NEORV32 RISC-V Processor, https://github.com/stnolting/neorv32                            #
-- # Copyright (c) 2024, Stephan Nolting. All rights reserved.                                     #
-- #                                                                                               #
-- # Redistribution and use in source and binary forms, with or without modification, are          #
-- # permitted provided that the following conditions are met:                                     #
-- #                                                                                               #
-- # 1. Redistributions of source code must retain the above copyright notice, this list of        #
-- #    conditions and the following disclaimer.                                                   #
-- #                                                                                               #
-- # 2. Redistributions in binary form must reproduce the above copyright notice, this list of     #
-- #    conditions and the following disclaimer in the documentation and/or other materials        #
-- #    provided with the distribution.                                                            #
-- #                                                                                               #
-- # 3. Neither the name of the copyright holder nor the names of its contributors may be used to  #
-- #    endorse or promote products derived from this software without specific prior written      #
-- #    permission.                                                                                #
-- #                                                                                               #
-- # THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS" AND ANY EXPRESS   #
-- # OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED WARRANTIES OF               #
-- # MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE    #
-- # COPYRIGHT HOLDER OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL,     #
-- # EXEMPLARY, OR CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE #
-- # GOODS OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER CAUSED    #
-- # AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT (INCLUDING     #
-- # NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED  #
-- # OF THE POSSIBILITY OF SUCH DAMAGE.                                                            #
-- #################################################################################################

library ieee;
use ieee.std_logic_1164.all;

library neorv32;
use neorv32.neorv32_package.all; -- the processor

library work;
use work.all; -- this module

library iCE40UP;
use iCE40UP.components.all; -- for device primitives

entity icebreaker_top is
  port ( -- add ports as required
    -- on-board USB-UART bridge --
    uart_txd_o  : out std_ulogic;
    uart_rxd_i  : in  std_ulogic;
    -- on-board SPI flash --
    flash_sck_o : out std_ulogic;
    flash_sdo_o : out std_ulogic;
    flash_sdi_i : in  std_ulogic;
    flash_csn_o : out std_ulogic;
    -- on-board LEDs --
    led_gr_o    : out std_ulogic; -- low-active green LED
    led_rd_o    : out std_ulogic; -- low-active red LED
    -- on-board user button --
    button_i    : in  std_ulogic  -- low-active reset button
  );
end icebreaker_top;

architecture icebreaker_top_rtl of icebreaker_top is

  -- configuration --
  constant f_clock_c : natural := 24000000; -- PLL output clock frequency in Hz

  -- on-chip oscillator --
  signal hf_osc_clk : std_logic;

  -- PLL (macro generated by radiant) --
  component system_pll
  port (
    ref_clk_i   : in  std_logic;
    rst_n_i     : in  std_logic;
    lock_o      : out std_logic;
    outcore_o   : out std_logic;
    outglobal_o : out std_logic
  );
  end component;
  --
  signal pll_rstn : std_logic;
  signal pll_lock : std_logic;
  signal pll_clk  : std_logic;

  -- CPU --
  signal cpu_clk  : std_ulogic;
  signal cpu_rstn : std_ulogic;

  -- internal IO connection --
  signal io_spi_sck : std_ulogic;
  signal io_spi_sdi : std_ulogic;
  signal io_spi_sdo : std_ulogic;
  signal io_spi_csn : std_ulogic_vector(7 downto 0);
  signal io_gpio_o  : std_ulogic_vector(63 downto 0);

begin

  -- On-Chip HF Oscillator (device primitive) -----------------------------------------------
  -- -------------------------------------------------------------------------------------------
  -- Clock divider selection: 0b00 = 48 MHz, 0b01 = 24 MHz, 0b10 = 12 MHz, 0b11 = 6 MHz
  HSOSC_inst : HSOSC
  generic map (
    CLKHF_DIV => "0b10" -- 12 MHz
  )
  port map (
    CLKHFPU => '1',
    CLKHFEN => '1',
    CLKHF   => hf_osc_clk
  );


  -- System PLL (macro generated as Lattice Radiant IP) -------------------------------------
  -- -------------------------------------------------------------------------------------------
  system_pll_inst: system_pll
  port map (
    ref_clk_i   => hf_osc_clk,
    rst_n_i     => pll_rstn,
    lock_o      => pll_lock,
    outcore_o   => open,
    outglobal_o => pll_clk
  );

  pll_rstn <= std_logic(button_i); -- reset PLL (and the whole system) via user button
  cpu_clk  <= std_ulogic(pll_clk);
  cpu_rstn <= std_ulogic(pll_lock);


  -- The Core of the Problem ----------------------------------------------------------------
  -- -------------------------------------------------------------------------------------------
  neorv32_inst: neorv32_top
  generic map ( -- add configuration options as required
    -- General --
    CLOCK_FREQUENCY   => f_clock_c, -- clock frequency of clk_i in Hz
    INT_BOOTLOADER_EN => true,      -- boot configuration: true = boot explicit bootloader; false = boot from int/ext (I)MEM

    -- RISC-V CPU Extensions --
    RISCV_ISA_A       => true,      -- implement atomic memory operations extension?
    RISCV_ISA_M       => true,      -- implement mul/div extension?
    RISCV_ISA_U       => true,      -- implement user mode extension?
    RISCV_ISA_Zicntr  => true,      -- implement base counters?
    RISCV_ISA_Zicond  => true,      -- implement integer conditional operations?

    -- Internal Instruction memory (IMEM) --
    MEM_INT_IMEM_EN   => true,      -- implement processor-internal instruction memory
    MEM_INT_IMEM_SIZE => 64*1024,   -- size of processor-internal instruction memory in bytes

    -- Internal Data memory (DMEM) --
    MEM_INT_DMEM_EN   => true,      -- implement processor-internal data memory
    MEM_INT_DMEM_SIZE => 64*1024,   -- size of processor-internal data memory in bytes

    -- Processor peripherals --
    IO_GPIO_NUM       => 32,        -- number of GPIO input/output pairs (0..64)
    IO_MTIME_EN       => true,      -- implement machine system timer (MTIME)?
    IO_UART0_EN       => true,      -- implement primary universal asynchronous receiver/transmitter (UART0)?
    IO_UART0_RX_FIFO  => 64,        -- RX fifo depth, has to be a power of two, min 1
    IO_UART0_TX_FIFO  => 64,        -- TX fifo depth, has to be a power of two, min 1
    IO_SPI_EN         => true,      -- implement serial peripheral interface (SPI)?
    IO_SPI_FIFO       => 1          -- SPI RTX fifo depth, has to be a power of two, min 1
  )
  port map ( -- add ports as required
    -- Global control --
    clk_i       => cpu_clk,
    rstn_i      => cpu_rstn,

    -- GPIO (available if IO_GPIO_NUM > 0) --
    gpio_o      => io_gpio_o,
    gpio_i      => (others => '0'),

    -- primary UART0 (available if IO_UART0_EN = true) --
    uart0_txd_o => uart_txd_o,
    uart0_rxd_i => uart_rxd_i,

    -- SPI (available if IO_SPI_EN = true) --
    spi_clk_o   => io_spi_sck,
    spi_dat_o   => io_spi_sdo,
    spi_dat_i   => io_spi_sdi,
    spi_csn_o   => io_spi_csn
  );


  -- IO Connection --------------------------------------------------------------------------
  -- -------------------------------------------------------------------------------------------

  -- on-board LEDs --
  led_gr_o <= not io_gpio_o(0); -- low-active
  led_rd_o <= not io_gpio_o(1); -- low-active

  -- on-board SPI flash --
  flash_sck_o <= io_spi_sck;
  flash_sdo_o <= io_spi_sdo;
  flash_csn_o <= io_spi_csn(0);
  io_spi_sdi  <= flash_sdi_i;


end icebreaker_top_rtl;
